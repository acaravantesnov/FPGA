--=================================================================================================
-- Title       : Comparator
-- File        : comparator_rtl.vhd
-- Description : Comparator entity for both the lfsr_seed_instance in lfsr sub-PUF, and for main
--               comparator.
--               As soon as the component stops receiving an active reset signal (either through
--               reset_n or aux_reset_n), from the first clk rising edge it starts counting RO clk
--               pulses. At the same time, an additional timer increments with the main clk of the
--               system. The g_timer_eoc indicates the component when to stop incrementing the
--               timer, and compare the number of pulses stored in each consecutive pair of RO clk
--               counters. This generates a value of width g_input_wdith / 2.
-- Generics    : g_input_width      -> Number of RO clks to compare.
--               g_timer_eoc        -> Final value of the timer counter. Value at which RO counters
--                                     are compared to generate the output.
--               g_reset_polarity   -> Active high ('1') or active low ('0') rest for both reset_n
--                                     and aux_reset_n.
-- Author      : Alberto Caravantes Arranz
-- Date        : 06/04/2025
-- Version     : 1.0
--=================================================================================================

-- Revision History:
-- Version 1.0 - Initial version

library ieee;
use ieee.std_logic_1164.all;

entity comparator is
    generic(
        g_input_width   : natural := 10;
        g_timer_eoc     : natural := 100E3;
        g_reset_polarity: std_logic := '0'
    );
    port(
        clk                 : in std_logic;
        aux_reset_n         : in std_logic;
        aux_2_reset_n       : in std_logic;
        reset_n             : in std_logic; -- Resets Counters and Timer, generated by FSM in lfsr_seed_inst, by input in comparator_inst
        RO_clks             : in std_logic_vector(g_input_width - 1 downto 0);
        comparison_result   : out std_logic_vector((g_input_width / 2) - 1 downto 0);
        value_ready         : out std_logic
    );
end entity comparator;

architecture rtl of comparator is

    constant c_output_width: natural := (g_input_width / 2);

    type t_natural_array is array (natural range <>) of natural;
    signal counter_i: t_natural_array(g_input_width - 1 downto 0);

    signal timer_i: natural range 0 to g_timer_eoc;
    signal eoc_i: std_logic;

    signal comparison_result_i: std_logic_vector(c_output_width - 1 downto 0);
    signal flag: std_logic;

begin

    GEN_COUNTERS: for i in 0 to g_input_width - 1 generate
        process(reset_n, aux_reset_n, aux_2_reset_n, RO_clks(i))
        begin
            if ((reset_n = g_reset_polarity) or (aux_reset_n = g_reset_polarity) or (aux_2_reset_n = g_reset_polarity))then
                counter_i(i) <= 0;
            elsif (rising_edge(RO_clks(i))) then
                if (eoc_i = '0') then
                    counter_i(i) <= counter_i(i) + 1;
                end if;
            end if;
        end process;
    end generate GEN_COUNTERS;

    PROC_TIMER: process(reset_n, aux_reset_n, aux_2_reset_n, clk)
    begin
        if ((reset_n = g_reset_polarity) or (aux_reset_n = g_reset_polarity) or (aux_2_reset_n = g_reset_polarity)) then
            timer_i <= 0;
            eoc_i <= '0';
        elsif (rising_edge(clk)) then
            if (timer_i = g_timer_eoc) then
                eoc_i <= '1';
            else
                timer_i <= timer_i + 1;
            end if;
        end if;
    end process PROC_TIMER;

    PROC_COMPARATOR: process(reset_n, aux_reset_n, aux_2_reset_n, clk)
    begin
        if ((reset_n = g_reset_polarity) or (aux_reset_n = g_reset_polarity) or (aux_2_reset_n = g_reset_polarity)) then
            comparison_result_i <= (others => '0');
        elsif (rising_edge(clk)) then
            if (eoc_i = '1') then
                for i in 0 to c_output_width - 1 loop
                    if (2 * i + 1 < g_input_width) and (counter_i(2 * i) > counter_i(2 * i + 1)) then
                        comparison_result_i(i) <= '1';
                    else
                        comparison_result_i(i) <= '0';
                    end if;
                end loop;
            end if;
        end if;
    end process PROC_COMPARATOR;

    comparison_result <= comparison_result_i;

    -- value_ready set to '1' one clock cycle after eoc to make sure value is readable
    -- (combinational comparison has had enough time to be done).
    PROC_VALUE_READY: process(reset_n, aux_reset_n, aux_2_reset_n, clk)
    begin
        if ((reset_n = g_reset_polarity) or (aux_reset_n = g_reset_polarity) or (aux_2_reset_n = g_reset_polarity)) then
            value_ready <= '0';
            flag <= '0';
        elsif (rising_edge(clk)) then
            if ((eoc_i = '1') and (flag = '0')) then
                value_ready <= '1';
                flag <= '1';
            else
                value_ready <= '0';
                -- Not updating flag to '0' to avoid a loop of pulses inm value_ready,
                -- just a single pulse even if eoc remains high.
            end if;
        end if;
    end process PROC_VALUE_READY;

end architecture rtl;
